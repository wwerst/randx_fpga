----------------------------------------
--! @file
--! @brief Template brief statement
--! @author Will Werst
--! @date   May 2021
----------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Common;


entity HashEngineTB is
end HashEngineTB;

architecture behavioral of HashEngineTB is
begin
end architecture behavioral;
